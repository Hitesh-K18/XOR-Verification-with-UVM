interface xor_interface(input logic clock);
  logic A,B,C;
endinterface